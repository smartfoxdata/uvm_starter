interface starter_if;
   logic clk;
   logic rst;
   logic [7:0] data;
   logic valid;
endinterface // starter_if
