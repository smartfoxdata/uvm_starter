`include "starter_if.sv"

package starter_pkg;

   import uvm_pkg::*;

`include "uvm_macros.svh"

`include "starter_txn.sv"
`include "starter_sqr.sv"
`include "starter_drv.sv"
`include "starter_mon.sv"
`include "starter_agt.sv"
`include "starter_env.sv"
`include "starter_seq_lib.sv"

endpackage // starter_pkg

